--
-- @author Peter Tisovcik <xtisov00@fit.vutbr.cz
--

library ieee;
use ieee.std_logic_1164.all;
library ieee;
use ieee.std_logic_1164.all;
-- ----------------------------------------------------------------------------
--                        Entity declaration
-- ----------------------------------------------------------------------------
entity fsm is
port(
   CLK         : in  std_logic;
   RESET       : in  std_logic;

   -- Input signals
   KEY         : in  std_logic_vector(15 downto 0);
   CNT_OF      : in  std_logic;

   -- Output signals
   FSM_CNT_CE  : out std_logic;
   FSM_MX_MEM  : out std_logic;
   FSM_MX_LCD  : out std_logic;
   FSM_LCD_WR  : out std_logic;
   FSM_LCD_CLR : out std_logic
);
end entity fsm;

-- ----------------------------------------------------------------------------
--                      Architecture declaration
-- ----------------------------------------------------------------------------
architecture behavioral of fsm is
   type t_state is (WAIT1, FAIL, TEST1, TEST2, TEST3, TEST4, TEST5, TEST6, TEST7,
   TEST8, TEST9, TEST10, TEST11, TEST12, TEST13, TEST14, TEST15, LAST_TEST,
   PRINT_MESSAGE_FAIL, PRINT_MESSAGE_SUCC, FINISH);
   signal present_state, next_state : t_state;

begin
-- -------------------------------------------------------
sync_logic : process(RESET, CLK)
begin
   if (RESET = '1') then
      present_state <= TEST1;
   elsif (CLK'event AND CLK = '1') then
      present_state <= next_state;
   end if;
end process sync_logic;

-- -------------------------------------------------------
next_state_logic : process(present_state, KEY, CNT_OF)
begin
   case (present_state) is
   -- - - - - - - - - - - - - - - - - - - - - - -
   when WAIT1 =>
      next_state <= TEST1;
   --
   when FAIL =>
      next_state <= FAIL;
      if (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      end if;

   -- TEST1 - 1
   when TEST1 =>
      next_state <= TEST1;
      if (KEY(1) = '1') then
         next_state <= TEST2;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST2 - 0
   when TEST2 =>
      next_state <= TEST2;
      if (KEY(0) = '1') then
         next_state <= TEST3;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST3 - 6
   when TEST3 =>
      next_state <= TEST3;
      if (KEY(6) = '1') then
         next_state <= TEST4;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST4 - 3
   when TEST4 =>
      next_state <= TEST4;
      if (KEY(3) = '1') then
         next_state <= TEST5;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST5 - 2 || 5
   when TEST5 =>
      next_state <= TEST5;
      if (KEY(2) = '1') then
         next_state <= TEST6;
	  elsif (KEY(5) = '1') then
	     next_state <= TEST11;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- prva varianta kodu
   -- TEST6 - 0
   when TEST6 =>
      next_state <= TEST6;
      if (KEY(0) = '1') then
         next_state <= TEST7;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST7 - 8
   when TEST7 =>
      next_state <= TEST7;
      if (KEY(8) = '1') then
         next_state <= TEST8;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST8 - 8
   when TEST8 =>
      next_state <= TEST8;
      if (KEY(8) = '1') then
         next_state <= TEST9;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST9 - 0
   when TEST9 =>
      next_state <= TEST9;
      if (KEY(0) = '1') then
         next_state <= TEST10;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST10 - 7
   when TEST10 =>
      next_state <= TEST10;
      if (KEY(7) = '1') then
         next_state <= LAST_TEST;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- pokracovanie druheho kodu
   -- TEST11 - 3
   when TEST11 =>
      next_state <= TEST11;
      if (KEY(3) = '1') then
         next_state <= TEST12;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST12 - 0
   when TEST12 =>
      next_state <= TEST12;
      if (KEY(0) = '1') then
         next_state <= TEST13;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST13 - 6
   when TEST13 =>
      next_state <= TEST13;
      if (KEY(6) = '1') then
         next_state <= TEST14;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST14 - 4
   when TEST14 =>
      next_state <= TEST14;
      if (KEY(4) = '1') then
         next_state <= TEST15;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- TEST15 - 2
   when TEST15 =>
      next_state <= TEST15;
      if (KEY(2) = '1') then
         next_state <= LAST_TEST;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_FAIL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- --------------------------------------------
   when LAST_TEST =>
      next_state <= LAST_TEST;
      if (KEY(15) = '1') then
         next_state <= PRINT_MESSAGE_SUCC;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;

   -- --------------------------------------------
   when PRINT_MESSAGE_SUCC =>
      next_state <= PRINT_MESSAGE_SUCC;
      if (CNT_OF = '1') then
         next_state <= FINISH;
      end if;

   -- --------------------------------------------
   when PRINT_MESSAGE_FAIL =>
      next_state <= PRINT_MESSAGE_FAIL;
      if (CNT_OF = '1') then
         next_state <= FINISH;
      end if;

   -- --------------------------------------------
   when FINISH =>
      next_state <= FINISH;
      if (KEY(15) = '1') then
         next_state <= TEST1;
      end if;

   -- --------------------------------------------
   when others =>
      next_state <= WAIT1;
   end case;
end process next_state_logic;

-- -------------------------------------------------------
output_logic : process(present_state, KEY)
begin
   FSM_CNT_CE     <= '0';
   FSM_MX_MEM     <= '0';
   FSM_MX_LCD     <= '0';
   FSM_LCD_WR     <= '0';
   FSM_LCD_CLR    <= '0';

   case (present_state) is
   -- - - - - - - - - - - - - - - - - - - - - - -
   when PRINT_MESSAGE_FAIL =>
      FSM_CNT_CE     <= '1';
      FSM_MX_LCD     <= '1';
      FSM_MX_MEM     <= '0';
      FSM_LCD_WR     <= '1';

   -- - - - - - - - - - - - - - - - - - - - - - -
   when PRINT_MESSAGE_SUCC =>
      FSM_CNT_CE     <= '1';
      FSM_MX_LCD     <= '1';
      FSM_MX_MEM     <= '1';
      FSM_LCD_WR     <= '1';

   -- - - - - - - - - - - - - - - - - - - - - - -
   when FINISH =>
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;

   -- - - - - - - - - - - - - - - - - - - - - - -
   when others =>
   if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
   end case;
end process output_logic;

end architecture behavioral;
